module fifo(clk,res,w_en,r_en,w_d,r_d);


endmodule
