class fifo_sbd;

        wr_tx w_t;
        rd_tx r_t;

        task run();
//            $display("FIFO_SBD is happening");
        endtask

endclass
