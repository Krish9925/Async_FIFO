class wr_cov;

        wr_tx tx;
        
        task run();
//            $display("WR_COV is happening");
        endtask

endclass
