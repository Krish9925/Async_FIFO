class rd_cov;

        rd_tx tx;
        
        task run();
//            $display("rd_COV is happening");
        endtask

endclass
