class rd_mon;

        rd_tx tx;

        task run();

//            $display("rd_MON is happening");

        endtask
endclass

