class rd_gen;

        rd_tx tx;

        task run();

//            $display("RD_TX is happening");

        endtask

endclass
