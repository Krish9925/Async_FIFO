class rd_bfm;

        rd_tx tx;

        task run();
//            $display("rd_BFM is happening");
        endtask

endclass
