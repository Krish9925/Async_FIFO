class wr_mon;

        wr_tx tx;

        task run();

//            $display("WR_MON is happening");

        endtask
endclass
